----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:05:56 01/08/2024 
-- Design Name: 
-- Module Name:    prueba_pmod - aprueba 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

use IEEE.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity prueba_pmod is
    Port ( 
			  clk : in std_logic;
			  boton : in std_logic;
			  col: out std_logic_vector(1 to 8);
			  filas : out std_logic_vector(1 to 8);
			  puntaje : out std_logic_vector(6 downto 0);
			  puntaje2: out std_logic_vector(6 downto 0);
			  mux : out std_logic_vector(3 downto 0));
end prueba_pmod;

architecture aprueba of prueba_pmod is

	signal clk_div : std_logic_vector(25 downto 0) := (OTHERS => '0');
	type Estados is (FRM_1, FRM_2, FRM_3, FRM_4, FRM_5, FRM_6, FRM_7, FRM_8, FRM_9, FRM_10, 
						  FRM_11, FRM_12, FRM_13, FRM_14, FRM_15, FRM_16, FRM_17, FRM_18, FRM_19, 
						  FRM_20, FRM_21, FRM_22, FRM_23, FRM_24, FRM_25, FRM_26, FRM_27, FRM_28, 
						  FRM_29, FRM_30, FRM_31, FRM_32, FRM_33, FRM_34, FRM_35, FRM_36, FRM_37, 
						  FRM_38, FRM_39, FRM_40, FRM_41, FRM_42, FRM_43, FRM_44, FRM_45, FRM_46, 
						  FRM_47, FRM_48, FRM_49, FRM_50, FRM_51, FRM_52, FRM_53, FRM_54, FRM_55, 
						  FRM_56, FRM_57, FRM_58, FRM_59, FRM_60, FRM_61, FRM_62, FRM_63, FRM_64, 
						  FRM_65, FRM_66, FRM_67, FRM_68, FRM_69, FRM_70, FRM_71, FRM_72, FRM_73, 
						  FRM_74, FRM_75, FRM_76, FRM_77, FRM_78, FRM_79, FRM_80, FRM_MUERTO0,
						  FRM_MUERTO1, FRM_MUERTO2, FRM_MUERTO3, FRM_MUERTO4, POR_10, POR_11, POR_12,
						  POR_13, POR_14, POR_15, POR_16, POR_17, POR_18, POR_19, POR_20, POR_21,
						  POR_22, POR_23, POR_24, POR_25, POR_26, POR_27, POR_28, POR_29, POR_30,
						  POR_31, POR_32, POR_33, POR_34, POR_35, POR_36, POR_37, POR_38, WIN_1, 
						  WIN_2, WIN_3, WIN_4, WIN_5, WIN_6, WIN_7, WIN_8, WIN_9, WIN_10, WIN_11, 
						  WIN_12, WIN_13, WIN_14, WIN_15, WIN_16, WIN_17, WIN_18, WIN_19, WIN_20, 
						  WIN_21, WIN_22, WIN_23, WIN_24, WIN_25, WIN_26, WIN_27, WIN_28, WIN_29,
						  WIN_30, WIN_31, WIN_32, WIN_33, WIN_34, WIN_35, WIN_36, WIN_37, WIN_38,
						  WIN_39, WIN_40, WIN_41, WIN_42, WIN_43, WIN_44, WIN_45);
	signal presente, siguiente : Estados;
	
	type Est_col is (C1, C2, C3, C4, C5, C6, C7, C8);
	signal Cpres, Csig : Est_col;
	
	type Est_fil is (F1, F2, F3, F4, F5, F6, F7, F8);
	signal Fpres, Fsig : Est_fil;
	
	type salto is (S0, S1, S2, S3, S4, S5, DEAD0, DEAD1, DEAD2, DEAD3, TROPHY0, TROPHY1, TROPHY2,
						TROPHY3, TROPHY4, TROPHY5, TROPHY6, TROPHY7, TROPHY8, FIN0, FIN1, FIN2, FIN3, 
						FIN4, FIN5);
	signal Spres, Ssig : salto;
	
	type matriz is array (1 to 8, 1 to 40) of std_logic;
	type tierra is array (1 to 8) of std_logic_vector(1 to 8);
	type seccion is array (1 to 8, 1 to 8) of std_logic;
	signal ventana : seccion;
	
	signal indice : integer range 1 to 8 := 1;
	signal score : integer range 0 to 10 := 0;
	
	constant Cuno 	  : std_logic_vector(1 to 8) := "10000000";											  
	constant Cdos 	  : std_logic_vector(1 to 8) := "01000000";
	constant Ctres   : std_logic_vector(1 to 8) := "00100000";
	constant Ccuatro : std_logic_vector(1 to 8) := "00010000";
	constant Ccinco  : std_logic_vector(1 to 8) := "00001000";
	constant Cseis   : std_logic_vector(1 to 8) := "00000100";
	constant Csiete  : std_logic_vector(1 to 8) := "00000010";
	constant Cocho   : std_logic_vector(1 to 8) := "00000001";									  
											  
	constant ESC_1 : seccion := (("11111001"),
								        ("11110000"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111110"),
								        ("00000000"));

	constant ESC_2 : seccion := (("11110011"),
								        ("11100001"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111101"),
								        ("00000000"));

	constant ESC_3 : seccion := (("11100111"),
								        ("11000011"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111011"),
								        ("00000000"));

	constant ESC_4 : seccion := (("11001111"),
								        ("10000111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11110111"),
								        ("00000000"));

	constant ESC_5 : seccion := (("10011111"),
								        ("00001111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11101111"),
								        ("00000000"));

	constant ESC_6 : seccion := (("00111111"),
								        ("00011110"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11011111"),
								        ("00000000"));

	constant ESC_7 : seccion := (("01111110"),
								        ("00111100"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("10111111"),
								        ("00000000"));

	constant ESC_8 : seccion := (("11111100"),
								        ("01111000"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("01111111"),
								        ("00000000"));

	constant ESC_9 : seccion := (("11111001"),
								        ("11110000"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_10 : seccion := (("11110011"),
								        ("11100001"),
								        ("11111111"),
								        ("11111111"),
								        ("11111110"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_11 : seccion := (("11100111"),
								        ("11000011"),
								        ("11111111"),
								        ("11111111"),
								        ("11111100"),
								        ("11111111"),
								        ("11111111"),
								        ("00000001"));

	constant ESC_12 : seccion := (("11001111"),
								        ("10000111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111000"),
								        ("11111111"),
								        ("11111111"),
								        ("00000010"));

	constant ESC_13 : seccion := (("10011111"),
								        ("00001111"),
								        ("11111111"),
								        ("11111111"),
								        ("11110000"),
								        ("11111111"),
								        ("11111111"),
								        ("00000100"));

	constant ESC_14 : seccion := (("00111111"),
								        ("00011110"),
								        ("11111111"),
								        ("11111111"),
								        ("11100000"),
								        ("11111111"),
								        ("11111111"),
								        ("00001000"));

	constant ESC_15 : seccion := (("01111110"),
								        ("00111100"),
								        ("11111111"),
								        ("11111111"),
								        ("11000001"),
								        ("11111111"),
								        ("11111111"),
								        ("00010000"));

	constant ESC_16 : seccion := (("11111100"),
								        ("01111000"),
								        ("11111111"),
								        ("11111111"),
								        ("10000011"),
								        ("11111111"),
								        ("11111111"),
								        ("00100000"));

	constant ESC_17 : seccion := (("11111001"),
								        ("11110000"),
								        ("11111111"),
								        ("11111111"),
								        ("00000111"),
								        ("11111111"),
								        ("11111111"),
								        ("01000000"));

	constant ESC_18 : seccion := (("11110011"),
								        ("11100001"),
								        ("11111111"),
								        ("11111111"),
								        ("00001111"),
								        ("11111111"),
								        ("11111111"),
								        ("10000000"));

	constant ESC_19 : seccion := (("11100111"),
								        ("11000011"),
								        ("11111111"),
								        ("11111111"),
								        ("00011111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_20 : seccion := (("11001111"),
								        ("10000111"),
								        ("11111111"),
								        ("11111111"),
								        ("00111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_21 : seccion := (("10011111"),
								        ("00001111"),
								        ("11111111"),
								        ("11111111"),
								        ("01111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_22 : seccion := (("00111111"),
								        ("00011110"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_23 : seccion := (("01111110"),
								        ("00111100"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_24 : seccion := (("11111100"),
								        ("01111000"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_25 : seccion := (("11111001"),
								        ("11110000"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_26 : seccion := (("11110011"),
								        ("11100001"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111110"),
								        ("00000000"));

	constant ESC_27 : seccion := (("11100111"),
								        ("11000011"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111101"),
								        ("00000000"));

	constant ESC_28 : seccion := (("11001111"),
								        ("10000111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111011"),
								        ("00000000"));

	constant ESC_29 : seccion := (("10011111"),
								        ("00001111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11110111"),
								        ("00000000"));

	constant ESC_30 : seccion := (("00111111"),
								        ("00011110"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11101111"),
								        ("00000000"));

	constant ESC_31 : seccion := (("01111110"),
								        ("00111100"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11011111"),
								        ("00000000"));

	constant ESC_32 : seccion := (("11111100"),
								        ("01111000"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("10111111"),
								        ("00000000"));

	constant ESC_33 : seccion := (("11111001"),
								        ("11110000"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("01111111"),
								        ("00000000"));

	constant ESC_34 : seccion := (("11110011"),
								        ("11100001"),
								        ("11111111"),
								        ("11111111"),
								        ("11111110"),
								        ("11111111"),
								        ("11111111"),
								        ("00000001"));

	constant ESC_35 : seccion := (("11100111"),
								        ("11000011"),
								        ("11111111"),
								        ("11111111"),
								        ("11111100"),
								        ("11111111"),
								        ("11111111"),
								        ("00000011"));

	constant ESC_36 : seccion := (("11001111"),
								        ("10000111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111000"),
								        ("11111111"),
								        ("11111111"),
								        ("00000111"));

	constant ESC_37 : seccion := (("10011111"),
								        ("00001111"),
								        ("11111111"),
								        ("11111111"),
								        ("11110000"),
								        ("11111111"),
								        ("11111111"),
								        ("00001111"));

	constant ESC_38 : seccion := (("00111111"),
								        ("00011110"),
								        ("11111111"),
								        ("11111111"),
								        ("11100000"),
								        ("11111111"),
								        ("11111111"),
								        ("00011111"));

	constant ESC_39 : seccion := (("01111110"),
								        ("00111100"),
								        ("11111111"),
								        ("11111111"),
								        ("11000000"),
								        ("11111111"),
								        ("11111111"),
								        ("00111111"));

	constant ESC_40 : seccion := (("11111100"),
								        ("01111000"),
								        ("11111111"),
								        ("11111111"),
								        ("10000000"),
								        ("11111111"),
								        ("11111111"),
								        ("01111111"));

	constant ESC_41 : seccion := (("11111001"),
								        ("11110000"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"));

	constant ESC_42 : seccion := (("11110011"),
								        ("11100001"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"));

	constant ESC_43 : seccion := (("11100111"),
								        ("11000011"),
								        ("11111111"),
								        ("11111111"),
								        ("00000001"),
								        ("11111111"),
								        ("11111111"),
								        ("11111110"));

	constant ESC_44 : seccion := (("11001111"),
								        ("10000111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000011"),
								        ("11111111"),
								        ("11111111"),
								        ("11111100"));

	constant ESC_45 : seccion := (("10011111"),
								        ("00001111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111000"));

	constant ESC_46 : seccion := (("00111111"),
								        ("00011110"),
								        ("11111111"),
								        ("11111111"),
								        ("00001111"),
								        ("11111111"),
								        ("11111111"),
								        ("11110000"));

	constant ESC_47 : seccion := (("01111110"),
								        ("00111100"),
								        ("11111111"),
								        ("11111111"),
								        ("00011111"),
								        ("11111111"),
								        ("11111111"),
								        ("11100000"));

	constant ESC_48 : seccion := (("11111100"),
								        ("01111000"),
								        ("11111111"),
								        ("11111111"),
								        ("00111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11000000"));

	constant ESC_49 : seccion := (("11111001"),
								        ("11110000"),
								        ("11111111"),
								        ("11111111"),
								        ("01111111"),
								        ("11111111"),
								        ("11111111"),
								        ("10000000"));

	constant ESC_50 : seccion := (("11110011"),
								        ("11100001"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_51 : seccion := (("11100111"),
								        ("11000011"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_52 : seccion := (("11001111"),
								        ("10000111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_53 : seccion := (("10011111"),
								        ("00001111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_54 : seccion := (("00111111"),
								        ("00011110"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_55 : seccion := (("01111110"),
								        ("00111100"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_56 : seccion := (("11111100"),
								        ("01111000"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000001"));

	constant ESC_57 : seccion := (("11111001"),
								        ("11110000"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000010"));

	constant ESC_58 : seccion := (("11110011"),
								        ("11100001"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000100"));

	constant ESC_59 : seccion := (("11100111"),
								        ("11000011"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00001000"));

	constant ESC_60 : seccion := (("11001111"),
								        ("10000111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00010000"));

	constant ESC_61 : seccion := (("10011111"),
								        ("00001111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00100000"));

	constant ESC_62 : seccion := (("00111111"),
								        ("00011111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("01000000"));

	constant ESC_63 : seccion := (("01111111"),
								        ("00111110"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("10000000"));

	constant ESC_64 : seccion := (("11111110"),
								        ("01111100"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000001"));

	constant ESC_65 : seccion := (("11111100"),
								        ("11111000"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000010"));

	constant ESC_66 : seccion := (("11111001"),
								        ("11110000"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111110"),
								        ("00000100"));

	constant ESC_67 : seccion := (("11110011"),
								        ("11100001"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111101"),
								        ("00001000"));

	constant ESC_68 : seccion := (("11100111"),
								        ("11000011"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111011"),
								        ("00010000"));

	constant ESC_69 : seccion := (("11001111"),
								        ("10000111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11110111"),
								        ("00100000"));

	constant ESC_70 : seccion := (("10011111"),
								        ("00001110"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11101111"),
								        ("01000000"));

	constant ESC_71 : seccion := (("00111110"),
								        ("00011100"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11011111"),
								        ("10000000"));

	constant ESC_72 : seccion := (("01111100"),
								        ("00111000"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("10111111"),
								        ("00000000"));

	constant ESC_73 : seccion := (("11111001"),
								        ("01110000"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("01111111"),
								        ("00000000"));

	constant ESC_74 : seccion := (("11110011"),
								        ("11100001"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_75 : seccion := (("11100111"),
								        ("11000011"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_76 : seccion := (("11001111"),
								        ("10000111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_77 : seccion := (("10011111"),
								        ("00001111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_78 : seccion := (("00111111"),
								        ("00011110"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_79 : seccion := (("01111110"),
								        ("00111100"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant ESC_80 : seccion := (("11111100"),
								        ("01111000"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("11111111"),
								        ("00000000"));

	constant MUERTO0 : seccion := (("10000001"),
											 ("00000000"),
											 ("00000000"),
											 ("00100100"),
											 ("00000000"),
											 ("11000011"),
											 ("11000011"),
											 ("11111111"));

	constant MUERTO1 : seccion := (("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"));

	constant MUERTO2 : seccion := (("10000001"),
											 ("00000000"),
											 ("00000000"),
											 ("00100100"),
											 ("00000000"),
											 ("11000011"),
											 ("11000011"),
											 ("11111111"));

	constant MUERTO3 : seccion := (("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"));

	constant MUERTO4 : seccion := (("10000001"),
											 ("00000000"),
											 ("00000000"),
											 ("00100100"),
											 ("00000000"),
											 ("11000011"),
											 ("11000011"),
											 ("11111111"));

	constant PORT_10 : seccion := (("11110011"),
								         ("11100001"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant PORT_11 : seccion := (("11100111"),
								         ("11000011"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000001"));

	constant PORT_12 : seccion := (("11001111"),
								         ("10000111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000010"));

	constant PORT_13 : seccion := (("10011111"),
								         ("00001111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000100"));

	constant PORT_14 : seccion := (("00111111"),
								         ("00011110"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00001000"));

	constant PORT_15 : seccion := (("01111110"),
								         ("00111100"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00010000"));

	constant PORT_16 : seccion := (("11111100"),
								         ("01111000"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00100000"));

	constant PORT_17 : seccion := (("11111001"),
								         ("11110000"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("01000000"));

	constant PORT_18 : seccion := (("11110011"),
								         ("11100001"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("10000000"));

	constant PORT_19 : seccion := (("11100111"),
								         ("11000011"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant PORT_20 : seccion := (("11001111"),
								         ("10000111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant PORT_21 : seccion := (("10011111"),
								         ("00001111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant PORT_22 : seccion := (("00111111"),
								         ("00011111"),
								         ("11111111"),
								         ("11111110"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant PORT_23 : seccion := (("01111111"),
								         ("00111111"),
								         ("11111110"),
								         ("11111100"),
								         ("11111110"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant PORT_24 : seccion := (("11111111"),
								         ("01111111"),
								         ("11111101"),
								         ("11111000"),
								         ("11111101"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant PORT_25 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111011"),
								         ("11110001"),
								         ("11111011"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant PORT_26 : seccion := (("11111111"),
								         ("11111111"),
								         ("11110111"),
								         ("11100011"),
								         ("11110111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant PORT_27 : seccion := (("11111111"),
								         ("11111111"),
								         ("11101111"),
								         ("11000111"),
								         ("11101111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant PORT_28 : seccion := (("11111111"),
								         ("11111111"),
								         ("11011111"),
								         ("10001111"),
								         ("11011111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant PORT_29 : seccion := (("11111111"),
								         ("11111111"),
								         ("10111111"),
								         ("00011111"),
								         ("10111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant PORT_30 : seccion := (("11111111"),
								         ("11111110"),
								         ("01111111"),
								         ("00111111"),
								         ("01111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant PORT_31 : seccion := (("11111110"),
								         ("11111100"),
								         ("11111111"),
								         ("01111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111110"),
								         ("00000000"));

	constant PORT_32 : seccion := (("11111100"),
								         ("11111000"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111101"),
								         ("00000000"));

	constant PORT_33 : seccion := (("11111001"),
								         ("11110000"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111011"),
								         ("00000000"));

	constant PORT_34 : seccion := (("11110011"),
								         ("11100001"),
								         ("11111111"),
								         ("11111111"),
								         ("11111110"),
								         ("11111111"),
								         ("11110111"),
								         ("00000001"));

	constant PORT_35 : seccion := (("11100111"),
								         ("11000011"),
								         ("11111111"),
								         ("11111111"),
								         ("11111100"),
								         ("11111111"),
								         ("11101111"),
								         ("00000011"));

	constant PORT_36 : seccion := (("11001111"),
								         ("10000111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111000"),
								         ("11111111"),
								         ("11011111"),
								         ("00000111"));

	constant PORT_37 : seccion := (("10011111"),
								         ("00001111"),
								         ("11111111"),
								         ("11111111"),
								         ("11110000"),
								         ("11111111"),
								         ("10111111"),
								         ("00001111"));

	constant PORT_38 : seccion := (("00111111"),
								         ("00011110"),
								         ("11111111"),
								         ("11111111"),
								         ("11100000"),
								         ("11111111"),
								         ("01111111"),
								         ("00011111"));

	constant GANA_1 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant GANA_2 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant GANA_3 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant GANA_4 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant GANA_5 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant GANA_6 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111110"),
								         ("00000000"));

	constant GANA_7 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111100"),
								         ("00000000"));

	constant GANA_8 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111110"),
								         ("11111000"),
								         ("00000000"));

	constant GANA_9 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111100"),
								         ("11110000"),
								         ("00000000"));

	constant GANA_10 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111110"),
								         ("11111000"),
								         ("11100000"),
								         ("00000000"));

	constant GANA_11 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111100"),
								         ("11110000"),
								         ("11000000"),
								         ("00000000"));

	constant GANA_12 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111000"),
								         ("11100000"),
								         ("10000000"),
								         ("00000000"));

	constant GANA_13 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11110000"),
								         ("11000000"),
								         ("00000000"),
								         ("00000000"));

	constant GANA_14 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11100000"),
								         ("10000000"),
								         ("00000000"),
								         ("00000000"));

	constant GANA_15 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11000000"),
								         ("00000000"),
								         ("00000000"),
								         ("00000000"));

	constant GANA_16 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("10000001"),
								         ("00000001"),
								         ("00000001"),
								         ("00000000"));

	constant GANA_17 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000011"),
								         ("00000011"),
								         ("00000011"),
								         ("00000000"));

	constant GANA_18 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000111"),
								         ("00000111"),
								         ("00000111"),
								         ("00000000"));

	constant GANA_19 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00001111"),
								         ("00001111"),
								         ("00001111"),
								         ("00000000"));

	constant GANA_20 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00011111"),
								         ("00011111"),
								         ("00011111"),
								         ("00000000"));

	constant GANA_21 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00111111"),
								         ("00111111"),
								         ("00111111"),
								         ("00000000"));

	constant GANA_22 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("01111111"),
								         ("01111111"),
								         ("01111111"),
								         ("00000000"));

	constant GANA_23 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant GANA_24 : seccion := (("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant GANA_25 : seccion := (("11111111"),
								         ("11111110"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant GANA_26 : seccion := (("11111111"),
								         ("11111100"),
								         ("11111110"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("11111111"),
								         ("00000000"));

	constant GANA_27 : seccion := (("11111111"),
								         ("11111000"),
								         ("11111100"),
								         ("11111110"),
								         ("11111110"),
								         ("11111110"),
								         ("11111110"),
								         ("00000000"));

	constant GANA_28 : seccion := (("11111111"),
								         ("11110001"),
								         ("11111001"),
								         ("11111101"),
								         ("11111101"),
								         ("11111101"),
								         ("11111101"),
								         ("00000000"));

	constant GANA_29 : seccion := (("11111111"),
								         ("11100011"),
								         ("11110011"),
								         ("11111011"),
								         ("11111011"),
								         ("11111011"),
								         ("11111011"),
								         ("00000000"));

	constant GANA_30 : seccion := (("11111111"),
								         ("11000111"),
								         ("11100111"),
								         ("11110111"),
								         ("11110111"),
								         ("11110111"),
								         ("11110111"),
								         ("00000000"));

	constant GANA_31 : seccion := (("11111111"),
								         ("10001111"),
								         ("11001111"),
								         ("11101111"),
								         ("11101111"),
								         ("11101111"),
								         ("11101111"),
								         ("00000000"));

	constant GANA_32 : seccion := (("11111111"),
								         ("00011111"),
								         ("10011111"),
								         ("11011111"),
								         ("11011111"),
								         ("11011111"),
								         ("11011111"),
								         ("00000000"));

	constant GANA_33 : seccion := (("11111111"),
								         ("00011111"),
								         ("10011111"),
								         ("11011111"),
								         ("11011111"),
								         ("11011111"),
								         ("11011111"),
								         ("00000000"));

	constant GANA_34 : seccion := (("11111111"),
								         ("00011111"),
								         ("10011111"),
								         ("11011111"),
								         ("11011111"),
								         ("11011111"),
								         ("11011111"),
								         ("00000000"));

	constant GANA_35 : seccion := (("11111111"),
								         ("00011111"),
								         ("10011111"),
								         ("11011111"),
								         ("11011111"),
								         ("11011111"),
								         ("11011111"),
								         ("00000000"));

	constant GANA_36 : seccion := (("11111111"),
								         ("00011111"),
								         ("10011111"),
								         ("11011111"),
								         ("11011111"),
								         ("11011111"),
								         ("11011111"),
								         ("00000000"));
											
	constant GANA_37 : seccion := (("11000011"),
											 ("00011000"),
											 ("01011010"),
											 ("10011001"),
											 ("11100111"),
											 ("11100111"),
											 ("11000011"),
											 ("11111111"));

											
	constant GANA_38 : seccion := (("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"));
											
	constant GANA_39 : seccion := (("11000011"),
											 ("00011000"),
											 ("01011010"),
											 ("10011001"),
											 ("11100111"),
											 ("11100111"),
											 ("11000011"),
											 ("11111111"));

											
	constant GANA_40 : seccion := (("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"),
											 ("11111111"));
											
	constant GANA_41 : seccion := (("11000011"),
											 ("00011000"),
											 ("01011010"),
											 ("10011001"),
											 ("11100111"),
											 ("11100111"),
											 ("11000011"),
											 ("11111111"));
											
	constant GANA_42 : seccion := (("11000011"),
											 ("00011000"),
											 ("01011010"),
											 ("10011001"),
											 ("11100111"),
											 ("11100111"),
											 ("11000011"),
											 ("11111111"));
											
	constant GANA_43 : seccion := (("11000011"),
											 ("00011000"),
											 ("01011010"),
											 ("10011001"),
											 ("11100111"),
											 ("11100111"),
											 ("11000011"),
											 ("11111111"));
											
	constant GANA_44 : seccion := (("11000011"),
											 ("00011000"),
											 ("01011010"),
											 ("10011001"),
											 ("11100111"),
											 ("11100111"),
											 ("11000011"),
											 ("11111111"));
											
	constant GANA_45 : seccion := (("11000011"),
											 ("00011000"),
											 ("01011010"),
											 ("10011001"),
											 ("11100111"),
											 ("11100111"),
											 ("11000011"),
											 ("11111111"));
			  
begin

	process (clk) begin
		if rising_edge(clk) then
			clk_div <= clk_div + '1';
		end if;
	end process;
	
	process (clk_div(15)) begin
		if rising_edge(clk_div(15)) then
			Cpres <= Csig;
			Fpres <= Fsig;
		end if;
	end process;

	process (Cpres) begin
		case (Cpres) is
			when C1 => col <= Cuno;
				Csig <= C2;
			when C2 => col <= Cdos;
				Csig <= C3;
			when C3 => col <= Ctres;
				Csig <= C4;
			when C4 => col <= Ccuatro;
				Csig <= C5;
			when C5 => col <= Ccinco;
				Csig <= C6;
			when C6 => col <= Cseis;
				Csig <= C7;
			when C7 => col <= Csiete;
				Csig <= C8;
			when C8 => col <= Cocho;
				Csig <= C1;
		end case;
		
		
		case (Fpres) is
			when F1 => 
				filas(1) <= ventana(1, 1);
				filas(2) <= ventana(2, 1);
				filas(3) <= ventana(3, 1);
				filas(4) <= ventana(4, 1);
				filas(5) <= ventana(5, 1);
				filas(6) <= ventana(6, 1);
				filas(7) <= ventana(7, 1);
				filas(8) <= ventana(8, 1);
				Fsig <= F2;
			when F2 => 
				filas(1) <= ventana(1, 2);
				filas(2) <= ventana(2, 2);
				filas(3) <= ventana(3, 2);
				filas(4) <= ventana(4, 2);
				filas(5) <= ventana(5, 2);
				filas(6) <= ventana(6, 2);
				filas(7) <= ventana(7, 2);
				filas(8) <= ventana(8, 2);
				Fsig <= F3;
			when F3 =>
				filas(1) <= ventana(1, 3);
				filas(2) <= ventana(2, 3);
				filas(3) <= ventana(3, 3);
				filas(4) <= ventana(4, 3);
				filas(5) <= ventana(5, 3);
				filas(6) <= ventana(6, 3);
				filas(7) <= ventana(7, 3);
				filas(8) <= ventana(8, 3);
				Fsig <= F4;
			when F4 =>
				filas(1) <= ventana(1, 4);
				filas(2) <= ventana(2, 4);
				filas(3) <= ventana(3, 4);
				filas(4) <= ventana(4, 4);
				filas(5) <= ventana(5, 4);
				filas(6) <= ventana(6, 4);
				filas(7) <= ventana(7, 4);
				filas(8) <= ventana(8, 4);
				Fsig <= F5;
			when F5 =>
				filas(1) <= ventana(1, 5);
				filas(2) <= ventana(2, 5);
				filas(3) <= ventana(3, 5);
				filas(4) <= ventana(4, 5);
				filas(5) <= ventana(5, 5);
				filas(6) <= ventana(6, 5);
				filas(7) <= ventana(7, 5);
				filas(8) <= ventana(8, 5);
				Fsig <= F6;
			when F6 => 
				filas(1) <= ventana(1, 6);
				filas(2) <= ventana(2, 6);
				filas(3) <= ventana(3, 6);
				filas(4) <= ventana(4, 6);
				filas(5) <= ventana(5, 6);
				filas(6) <= ventana(6, 6);
				filas(7) <= ventana(7, 6);
				filas(8) <= ventana(8, 6);
				Fsig <= F7;
			when F7 => 
				filas(1) <= ventana(1, 7);
				filas(2) <= ventana(2, 7);
				filas(3) <= ventana(3, 7);
				filas(4) <= ventana(4, 7);
				filas(5) <= ventana(5, 7);
				filas(6) <= ventana(6, 7);
				filas(7) <= ventana(7, 7);
				filas(8) <= ventana(8, 7);
				Fsig <= F8;
			when F8 =>
				filas(1) <= ventana(1, 8);
				filas(2) <= ventana(2, 8);
				filas(3) <= ventana(3, 8);
				filas(4) <= ventana(4, 8);
				filas(5) <= ventana(5, 8);
				filas(6) <= ventana(6, 8);
				filas(7) <= ventana(7, 8);
				filas(8) <= ventana(8, 8);
				Fsig <= F1;
		end case;
	end process;
	
	process (clk_div(24)) begin
		if rising_edge(clk_div(24)) then
			if presente = WIN_45 then
				score <= 0;
			end if;
			presente <= siguiente;
			Spres <= Ssig;
			if	Spres = S0 then				
				if	score > 8 then
					presente <= WIN_1;
				end if;
			end if;
			if Spres = S5 then
				if ventana(7, 1) = '0' then
					score <= score + 1;
				end if;
			elsif Spres = S0 then -- MORIR
				if (presente = FRM_8) or (presente = FRM_33) or (presente = FRM_73) or -- ENEMIGOS FRM
					-- HUECOS FRM
					(presente = FRM_18) or (presente = FRM_41) or (presente = FRM_42) or
					(presente = FRM_43) or (presente = FRM_63) or (presente = FRM_71) or
					(presente = POR_18) or (presente = POR_38) then -- ENEMIGO y HUECO POR
					score <= 0;
					presente <= FRM_MUERTO0;
				end if;
			end if;
		end if;
	end process;
	
	process (presente) begin
		case (presente) is
			when FRM_1 => ventana <= ESC_1;
				siguiente <= FRM_2;
			when FRM_2 => ventana <= ESC_2;
				siguiente <= FRM_3;
			when FRM_3 => ventana <= ESC_3;
				siguiente <= FRM_4;
			when FRM_4 => ventana <= ESC_4;
				siguiente <= FRM_5;
			when FRM_5 => ventana <= ESC_5;
				siguiente <= FRM_6;
			when FRM_6 => ventana <= ESC_6;
				siguiente <= FRM_7;
			when FRM_7 => ventana <= ESC_7;
				siguiente <= FRM_8;
			when FRM_8 => ventana <= ESC_8;
				siguiente <= FRM_9;
			when FRM_9 => ventana <= ESC_9;
				if score > 4 then
					siguiente <= POR_10;
				else
					siguiente <= FRM_10;
				end if;
			when FRM_10 => ventana <= ESC_10;
				siguiente <= FRM_11;
			when FRM_11 => ventana <= ESC_11;
				siguiente <= FRM_12;
			when FRM_12 => ventana <= ESC_12;
				siguiente <= FRM_13;
			when FRM_13 => ventana <= ESC_13;
				siguiente <= FRM_14;
			when FRM_14 => ventana <= ESC_14;
				siguiente <= FRM_15;
			when FRM_15 => ventana <= ESC_15;
				siguiente <= FRM_16;
			when FRM_16 => ventana <= ESC_16;
				siguiente <= FRM_17;
			when FRM_17 => ventana <= ESC_17;
				siguiente <= FRM_18;
			when FRM_18 => ventana <= ESC_18;
				siguiente <= FRM_19;
			when FRM_19 => ventana <= ESC_19;
				siguiente <= FRM_20;
			when FRM_20 => ventana <= ESC_20;
				siguiente <= FRM_21;
			when FRM_21 => ventana <= ESC_21;
				siguiente <= FRM_22;
			when FRM_22 => ventana <= ESC_22;
				siguiente <= FRM_23;
			when FRM_23 => ventana <= ESC_23;
				siguiente <= FRM_24;
			when FRM_24 => ventana <= ESC_24;
				siguiente <= FRM_25;
			when FRM_25 => ventana <= ESC_25;
				siguiente <= FRM_26;
			when FRM_26 => ventana <= ESC_26;
				siguiente <= FRM_27;
			when FRM_27 => ventana <= ESC_27;
				siguiente <= FRM_28;
			when FRM_28 => ventana <= ESC_28;
				siguiente <= FRM_29;
			when FRM_29 => ventana <= ESC_29;
				siguiente <= FRM_30;
			when FRM_30 => ventana <= ESC_30;
				siguiente <= FRM_31;
			when FRM_31 => ventana <= ESC_31;
				siguiente <= FRM_32;
			when FRM_32 => ventana <= ESC_32;
				siguiente <= FRM_33;
			when FRM_33 => ventana <= ESC_33;
				siguiente <= FRM_34;
			when FRM_34 => ventana <= ESC_34;
				siguiente <= FRM_35;
			when FRM_35 => ventana <= ESC_35;
				siguiente <= FRM_36;
			when FRM_36 => ventana <= ESC_36;
				siguiente <= FRM_37;
			when FRM_37 => ventana <= ESC_37;
				siguiente <= FRM_38;
			when FRM_38 => ventana <= ESC_38;
				siguiente <= FRM_39;
			when FRM_39 => ventana <= ESC_39;
				siguiente <= FRM_40;
			when FRM_40 => ventana <= ESC_40;
				siguiente <= FRM_41;
			when FRM_41 => ventana <= ESC_41;
				siguiente <= FRM_42;
			when FRM_42 => ventana <= ESC_42;
				siguiente <= FRM_43;
			when FRM_43 => ventana <= ESC_43;
				siguiente <= FRM_44;
			when FRM_44 => ventana <= ESC_44;
				siguiente <= FRM_45;
			when FRM_45 => ventana <= ESC_45;
				siguiente <= FRM_46;
			when FRM_46 => ventana <= ESC_46;
				siguiente <= FRM_47;
			when FRM_47 => ventana <= ESC_47;
				siguiente <= FRM_48;
			when FRM_48 => ventana <= ESC_48;
				siguiente <= FRM_49;
			when FRM_49 => ventana <= ESC_49;
				siguiente <= FRM_50;
			when FRM_50 => ventana <= ESC_50;
				siguiente <= FRM_51;
			when FRM_51 => ventana <= ESC_51;
				siguiente <= FRM_52;
			when FRM_52 => ventana <= ESC_52;
				siguiente <= FRM_53;
			when FRM_53 => ventana <= ESC_53;
				siguiente <= FRM_54;
			when FRM_54 => ventana <= ESC_54;
				siguiente <= FRM_55;
			when FRM_55 => ventana <= ESC_55;
				siguiente <= FRM_56;
			when FRM_56 => ventana <= ESC_56;
				siguiente <= FRM_57;
			when FRM_57 => ventana <= ESC_57;
				siguiente <= FRM_58;
			when FRM_58 => ventana <= ESC_58;
				siguiente <= FRM_59;
			when FRM_59 => ventana <= ESC_59;
				siguiente <= FRM_60;
			when FRM_60 => ventana <= ESC_60;
				siguiente <= FRM_61;
			when FRM_61 => ventana <= ESC_61;
				siguiente <= FRM_62;
			when FRM_62 => ventana <= ESC_62;
				siguiente <= FRM_63;
			when FRM_63 => ventana <= ESC_63;
				siguiente <= FRM_64;
			when FRM_64 => ventana <= ESC_64;
				siguiente <= FRM_65;
			when FRM_65 => ventana <= ESC_65;
				siguiente <= FRM_66;
			when FRM_66 => ventana <= ESC_66;
				siguiente <= FRM_67;
			when FRM_67 => ventana <= ESC_67;
				siguiente <= FRM_68;
			when FRM_68 => ventana <= ESC_68;
				siguiente <= FRM_69;
			when FRM_69 => ventana <= ESC_69;
				siguiente <= FRM_70;
			when FRM_70 => ventana <= ESC_70;
				siguiente <= FRM_71;
			when FRM_71 => ventana <= ESC_71;
				siguiente <= FRM_72;
			when FRM_72 => ventana <= ESC_72;
				siguiente <= FRM_73;
			when FRM_73 => ventana <= ESC_73;
				siguiente <= FRM_74;
			when FRM_74 => ventana <= ESC_74;
				siguiente <= FRM_75;
			when FRM_75 => ventana <= ESC_75;
				siguiente <= FRM_76;
			when FRM_76 => ventana <= ESC_76;
				siguiente <= FRM_77;
			when FRM_77 => ventana <= ESC_77;
				siguiente <= FRM_78;
			when FRM_78 => ventana <= ESC_78;
				siguiente <= FRM_79;
			when FRM_79 => ventana <= ESC_79;
				siguiente <= FRM_80;
			when FRM_80 => ventana <= ESC_80;
				siguiente <= FRM_1;
			when FRM_MUERTO0 => ventana <= MUERTO0;
				siguiente <= FRM_MUERTO1;
			when FRM_MUERTO1 => ventana <= MUERTO1;
				siguiente <= FRM_MUERTO2;
			when FRM_MUERTO2 => ventana <= MUERTO2;
				siguiente <= FRM_MUERTO3;
			when FRM_MUERTO3 => ventana <= MUERTO3;
				siguiente <= FRM_MUERTO4;
			when FRM_MUERTO4 => ventana <= MUERTO4;
				siguiente <= FRM_1;
			when POR_10 => ventana <= PORT_10;
				siguiente <= POR_11;
			when POR_11 => ventana <= PORT_11;
				siguiente <= POR_12;
			when POR_12 => ventana <= PORT_12;
				siguiente <= POR_13;
			when POR_13 => ventana <= PORT_13;
				siguiente <= POR_14;
			when POR_14 => ventana <= PORT_14;
				siguiente <= POR_15;
			when POR_15 => ventana <= PORT_15;
				siguiente <= POR_16;
			when POR_16 => ventana <= PORT_16;
				siguiente <= POR_17;
			when POR_17 => ventana <= PORT_17;
				siguiente <= POR_18;
			when POR_18 => ventana <= PORT_18;
				siguiente <= POR_19;
			when POR_19 => ventana <= PORT_19;
				siguiente <= POR_20;
			when POR_20 => ventana <= PORT_20;
				siguiente <= POR_21;
			when POR_21 => ventana <= PORT_21;
				siguiente <= POR_22;
			when POR_22 => ventana <= PORT_22;
				siguiente <= POR_23;
			when POR_23 => ventana <= PORT_23;
				siguiente <= POR_24;
			when POR_24 => ventana <= PORT_24;
				siguiente <= POR_25;
			when POR_25 => ventana <= PORT_25;
				siguiente <= POR_26;
			when POR_26 => ventana <= PORT_26;
				siguiente <= POR_27;
			when POR_27 => ventana <= PORT_27;
				siguiente <= POR_28;
			when POR_28 => ventana <= PORT_28;
				siguiente <= POR_29;
			when POR_29 => ventana <= PORT_29;
				if	Spres = S3 then
					siguiente <= WIN_1;
				else
					siguiente <= POR_30;
				end if;
			when POR_30 => ventana <= PORT_30;
				if	Spres = S3 then
					siguiente <= WIN_1;
				else
					siguiente <= POR_31;
				end if;
			when POR_31 => ventana <= PORT_31;
				if	Spres = S3 then
					siguiente <= WIN_1;
				else
					siguiente <= POR_32;
				end if;
			when POR_32 => ventana <= PORT_32;
				siguiente <= POR_33;
			when POR_33 => ventana <= PORT_33;
				siguiente <= POR_34;
			when POR_34 => ventana <= PORT_34;
				siguiente <= POR_35;
			when POR_35 => ventana <= PORT_35;
				siguiente <= POR_36;
			when POR_36 => ventana <= PORT_36;
				siguiente <= POR_37;
			when POR_37 => ventana <= PORT_37;
				siguiente <= POR_38;
			when POR_38 => ventana <= PORT_38;
				siguiente <= FRM_39;
			when WIN_1 => ventana <= GANA_1;
				siguiente <= WIN_2;
			when WIN_2 => ventana <= GANA_2;
				siguiente <= WIN_3;
			when WIN_3 => ventana <= GANA_3;
				siguiente <= WIN_4;
			when WIN_4 => ventana <= GANA_4;
				siguiente <= WIN_5;
			when WIN_5 => ventana <= GANA_5;
				siguiente <= WIN_6;
			when WIN_6 => ventana <= GANA_6;
				siguiente <= WIN_7;
			when WIN_7 => ventana <= GANA_7;
				siguiente <= WIN_8;
			when WIN_8 => ventana <= GANA_8;
				siguiente <= WIN_9;
			when WIN_9 => ventana <= GANA_9;
				siguiente <= WIN_10;
			when WIN_10 => ventana <= GANA_10;
				siguiente <= WIN_11;
			when WIN_11 => ventana <= GANA_11;
				siguiente <= WIN_12;
			when WIN_12 => ventana <= GANA_12;
				siguiente <= WIN_13;
			when WIN_13 => ventana <= GANA_13;
				siguiente <= WIN_14;
			when WIN_14 => ventana <= GANA_14;
				siguiente <= WIN_15;
			when WIN_15 => ventana <= GANA_15;
				siguiente <= WIN_16;
			when WIN_16 => ventana <= GANA_16;
				siguiente <= WIN_17;
			when WIN_17 => ventana <= GANA_17;
				siguiente <= WIN_18;
			when WIN_18 => ventana <= GANA_18;
				siguiente <= WIN_19;
			when WIN_19 => ventana <= GANA_19;
				siguiente <= WIN_20;
			when WIN_20 => ventana <= GANA_20;
				siguiente <= WIN_21;
			when WIN_21 => ventana <= GANA_21;
				siguiente <= WIN_22;
			when WIN_22 => ventana <= GANA_22;
				siguiente <= WIN_23;
			when WIN_23 => ventana <= GANA_23;
				siguiente <= WIN_24;
			when WIN_24 => ventana <= GANA_24;
				siguiente <= WIN_25;
			when WIN_25 => ventana <= GANA_25;
				siguiente <= WIN_26;
			when WIN_26 => ventana <= GANA_26;
				siguiente <= WIN_27;
			when WIN_27 => ventana <= GANA_27;
				siguiente <= WIN_28;
			when WIN_28 => ventana <= GANA_28;
				siguiente <= WIN_29;
			when WIN_29 => ventana <= GANA_29;
				siguiente <= WIN_30;
			when WIN_30 => ventana <= GANA_30;
				siguiente <= WIN_31;
			when WIN_31 => ventana <= GANA_31;
				siguiente <= WIN_32;
			when WIN_32 => ventana <= GANA_32;
				siguiente <= WIN_33;
			when WIN_33 => ventana <= GANA_33;
				siguiente <= WIN_34;
			when WIN_34 => ventana <= GANA_34;
				siguiente <= WIN_35;
			when WIN_35 => ventana <= GANA_35;
				siguiente <= WIN_36;
			when WIN_36 => ventana <= GANA_36;
				siguiente <= WIN_37;
			when WIN_37 => ventana <= GANA_37;
				siguiente <= WIN_38;
			when WIN_38 => ventana <= GANA_38;
				siguiente <= WIN_39;
			when WIN_39 => ventana <= GANA_39;
				siguiente <= WIN_40;
			when WIN_40 => ventana <= GANA_40;
				siguiente <= WIN_41;
			when WIN_41 => ventana <= GANA_41;
				siguiente <= WIN_42;
			when WIN_42 => ventana <= GANA_42;
				siguiente <= WIN_43;
			when WIN_43 => ventana <= GANA_43;
				siguiente <= WIN_44;
			when WIN_44 => ventana <= GANA_44;
				siguiente <= WIN_45;
			when WIN_45 => ventana <= GANA_45;
				siguiente <= FRM_1;
		end case;
		case (Spres) is
			when S0 =>
				if (presente = FRM_MUERTO0) then
					ventana(7, 1) <= '1';
					Ssig <= DEAD0;
				elsif (presente = WIN_1) or (presente = WIN_2) or (presente = WIN_3) or 
						(presente = WIN_4) or (presente = WIN_5) then
					ventana(7, 1) <= '0';
					Ssig <= FIN0;
				elsif boton = '1' then
					ventana(7, 1) <= '0';
					Ssig <= S1;
				else
					ventana(7, 1) <= '0';
					Ssig <= S0;
				end if;
			when S1 => ventana(6, 1) <= '0';
				Ssig <= S2;
			when S2 => ventana(5, 1) <= '0';
				Ssig <= S3;
			when S3 => ventana(4, 1) <= '0';
				if (presente = FRM_17) or (presente = FRM_18) or (presente = FRM_19) or 
					(presente = FRM_20) or (presente = FRM_21) or
					(presente = FRM_41) or (presente = FRM_42) or (presente = FRM_43) or 
					(presente = FRM_44) or (presente = FRM_45) or (presente = FRM_46) or 
					(presente = FRM_47) or (presente = FRM_48) or (presente = FRM_49) then
					Ssig <= S3;
				else
					Ssig <= S4;
				end if;
			when S4 => ventana(5, 1) <= '0';
				Ssig <= S5;
			when S5 => ventana(6, 1) <= '0';
				Ssig <= S0;
			when DEAD0 => ventana(7,1) <= '1';
				Ssig <= DEAD1;
			when DEAD1 => ventana(7,1) <= '1';
				Ssig <= DEAD2;
			when DEAD2 => ventana(7,1) <= '1';
				Ssig <= DEAD3;
			when DEAD3 => ventana(7,1) <= '1';
				Ssig <= S0;
			when FIN0 => ventana(7, 1) <= '0';
				if presente = WIN_11 then
					Ssig <= FIN1;
				elsif presente = WIN_36 then
					Ssig <= TROPHY0;
				else
					Ssig <= FIN0;
				end if;
			when FIN1 => ventana(6, 1) <= '0';
				if presente = WIN_13 then
					Ssig <= FIN2;
				else
					Ssig <= FIN1;
				end if;
			when FIN2 => ventana(5, 1) <= '0';
				if presente = WIN_15 then
					Ssig <= FIN3;
				else
					Ssig <= FIN2;
				end if;
			when FIN3 => ventana(4, 1) <= '0';
				if presente = WIN_23 then
					Ssig <= FIN4;
				else
					Ssig <= FIN3;
				end if;
			when FIN4 => ventana(5, 1) <= '0';
				Ssig <= FIN5;
			when FIN5 => ventana(6, 1) <= '0';
				Ssig <= FIN0;
			when TROPHY0 => ventana(7,1) <= '1';
				Ssig <= TROPHY1;
			when TROPHY1 => ventana(7,1) <= '1';
				Ssig <= TROPHY2;
			when TROPHY2 => ventana(7,1) <= '1';
				Ssig <= TROPHY3;
			when TROPHY3 => ventana(7,1) <= '1';
				Ssig <= TROPHY4;
			when TROPHY4 => ventana(7,1) <= '1';
				Ssig <= TROPHY5;
			when TROPHY5 => ventana(7,1) <= '1';
				Ssig <= TROPHY6;
			when TROPHY6 => ventana(7,1) <= '1';
				Ssig <= TROPHY7;
			when TROPHY7 => ventana(7,1) <= '1';
				Ssig <= TROPHY8;
			when TROPHY8 => ventana(7,1) <= '1';
				Ssig <= S0;
		end case;
	end process;
	
	process (score) begin
		case (score) is
			when 0 => puntaje <= "0000001";
				mux <= "1110";
			when 1 => puntaje <= "1001111";
				mux <= "1110";
			when 2 => puntaje <= "0010010";
				mux <= "1110";
			when 3 => puntaje <= "0000110";
				mux <= "1110";
			when 4 => puntaje <= "1001100";
				mux <= "1110";
			when 5 => puntaje <= "0100100";
				mux <= "1110";
			when 6 => puntaje <= "0100000";
				mux <= "1110";
			when 7 => puntaje <= "0001111";
				mux <= "1110";
			when 8 => puntaje <= "0000000";
				mux <= "1110";
			when 9 => puntaje <= "0000100";
				mux <= "1110";
			when others => puntaje <= "1111110";
				mux <= "1110";
		end case;
	end process;
	
end aprueba;

